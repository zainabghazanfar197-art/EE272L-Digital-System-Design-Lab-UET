module and_gate2 (
    input  logic A,
    input  logic B,
    output logic Y
);

    assign Y = A & B;

endmodule
